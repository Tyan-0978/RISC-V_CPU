// -----------------------------------------------------------------------------
// ALU top module
// -----------------------------------------------------------------------------

module alu (
    input  i_rst_n,
    input  i_clk,
    input  [?:0]  i_mode, // TODO
    input  [31:0] i_a,
    input  [31:0] i_b,
    output [31:0] o_result,
    output o_stall
);

// registers & wires -------------------------------------------------
// sub-module ports

// control signals

// sub-modules -------------------------------------------------------
// TODO

endmodule
