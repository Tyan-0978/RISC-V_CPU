// -----------------------------------------------------------------------------
// INT multiplication module
// -----------------------------------------------------------------------------

module int_mul (
    input  signed [31:0] i_a,
    input  signed [31:0] i_b,
    output signed [31:0] o_result
);

endmodule
