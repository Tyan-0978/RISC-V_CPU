module ecall (
    input 
    
    
    
    )


endmodule